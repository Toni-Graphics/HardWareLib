module main();
    initial begin
        $monitor("Write your code here");
    end
endmodule